// helen.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module helen (
		output wire        adc_sclk,                     //                   adc.sclk
		output wire        adc_cs_n,                     //                      .cs_n
		input  wire        adc_dout,                     //                      .dout
		output wire        adc_din,                      //                      .din
		input  wire        altpll_areset_conduit_export, // altpll_areset_conduit.export
		output wire        altpll_locked_conduit_export, // altpll_locked_conduit.export
		output wire        altpll_sdram_clk,             //          altpll_sdram.clk
		input  wire        clk_clk,                      //                   clk.clk
		output wire        flash_dclk,                   //                 flash.dclk
		output wire        flash_sce,                    //                      .sce
		output wire        flash_sdo,                    //                      .sdo
		input  wire        flash_data0,                  //                      .data0
		output wire [7:0]  ledg_export,                  //                  ledg.export
		input  wire        reset_reset_n,                //                 reset.reset_n
		output wire [12:0] sdram_wire_addr,              //            sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                //                      .ba
		output wire        sdram_wire_cas_n,             //                      .cas_n
		output wire        sdram_wire_cke,               //                      .cke
		output wire        sdram_wire_cs_n,              //                      .cs_n
		inout  wire [15:0] sdram_wire_dq,                //                      .dq
		output wire [1:0]  sdram_wire_dqm,               //                      .dqm
		output wire        sdram_wire_ras_n,             //                      .ras_n
		output wire        sdram_wire_we_n,              //                      .we_n
		input  wire        spi_MISO,                     //                   spi.MISO
		output wire        spi_MOSI,                     //                      .MOSI
		output wire        spi_SCLK,                     //                      .SCLK
		output wire        spi_SS_n,                     //                      .SS_n
		input  wire        uart_rxd,                     //                  uart.rxd
		output wire        uart_txd                      //                      .txd
	);

	wire         altpll_c0_clk;                                               // altpll:c0 -> [adc:clock, flash:clk, irq_mapper:clk, irq_mapper_001:clk, jtag_uart_0:clk, led:clk, mm_interconnect_0:altpll_c0_clk, nios_1:clk, nios_2:clk, onchip_1:clk, onchip_2:clk, rst_controller:clk, rst_controller_002:clk, rst_controller_003:clk, sdram:clk, spi_0:clk, sysid_qsys_1:clock, uart:clk]
	wire  [31:0] nios_1_data_master_readdata;                                 // mm_interconnect_0:nios_1_data_master_readdata -> nios_1:d_readdata
	wire         nios_1_data_master_waitrequest;                              // mm_interconnect_0:nios_1_data_master_waitrequest -> nios_1:d_waitrequest
	wire         nios_1_data_master_debugaccess;                              // nios_1:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios_1_data_master_debugaccess
	wire  [26:0] nios_1_data_master_address;                                  // nios_1:d_address -> mm_interconnect_0:nios_1_data_master_address
	wire   [3:0] nios_1_data_master_byteenable;                               // nios_1:d_byteenable -> mm_interconnect_0:nios_1_data_master_byteenable
	wire         nios_1_data_master_read;                                     // nios_1:d_read -> mm_interconnect_0:nios_1_data_master_read
	wire         nios_1_data_master_write;                                    // nios_1:d_write -> mm_interconnect_0:nios_1_data_master_write
	wire  [31:0] nios_1_data_master_writedata;                                // nios_1:d_writedata -> mm_interconnect_0:nios_1_data_master_writedata
	wire  [31:0] nios_2_data_master_readdata;                                 // mm_interconnect_0:nios_2_data_master_readdata -> nios_2:d_readdata
	wire         nios_2_data_master_waitrequest;                              // mm_interconnect_0:nios_2_data_master_waitrequest -> nios_2:d_waitrequest
	wire         nios_2_data_master_debugaccess;                              // nios_2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios_2_data_master_debugaccess
	wire  [26:0] nios_2_data_master_address;                                  // nios_2:d_address -> mm_interconnect_0:nios_2_data_master_address
	wire   [3:0] nios_2_data_master_byteenable;                               // nios_2:d_byteenable -> mm_interconnect_0:nios_2_data_master_byteenable
	wire         nios_2_data_master_read;                                     // nios_2:d_read -> mm_interconnect_0:nios_2_data_master_read
	wire         nios_2_data_master_write;                                    // nios_2:d_write -> mm_interconnect_0:nios_2_data_master_write
	wire  [31:0] nios_2_data_master_writedata;                                // nios_2:d_writedata -> mm_interconnect_0:nios_2_data_master_writedata
	wire  [31:0] nios_2_instruction_master_readdata;                          // mm_interconnect_0:nios_2_instruction_master_readdata -> nios_2:i_readdata
	wire         nios_2_instruction_master_waitrequest;                       // mm_interconnect_0:nios_2_instruction_master_waitrequest -> nios_2:i_waitrequest
	wire  [26:0] nios_2_instruction_master_address;                           // nios_2:i_address -> mm_interconnect_0:nios_2_instruction_master_address
	wire         nios_2_instruction_master_read;                              // nios_2:i_read -> mm_interconnect_0:nios_2_instruction_master_read
	wire  [31:0] nios_1_instruction_master_readdata;                          // mm_interconnect_0:nios_1_instruction_master_readdata -> nios_1:i_readdata
	wire         nios_1_instruction_master_waitrequest;                       // mm_interconnect_0:nios_1_instruction_master_waitrequest -> nios_1:i_waitrequest
	wire  [26:0] nios_1_instruction_master_address;                           // nios_1:i_address -> mm_interconnect_0:nios_1_instruction_master_address
	wire         nios_1_instruction_master_read;                              // nios_1:i_read -> mm_interconnect_0:nios_1_instruction_master_read
	wire  [31:0] mm_interconnect_0_adc_adc_slave_readdata;                    // adc:readdata -> mm_interconnect_0:adc_adc_slave_readdata
	wire         mm_interconnect_0_adc_adc_slave_waitrequest;                 // adc:waitrequest -> mm_interconnect_0:adc_adc_slave_waitrequest
	wire   [2:0] mm_interconnect_0_adc_adc_slave_address;                     // mm_interconnect_0:adc_adc_slave_address -> adc:address
	wire         mm_interconnect_0_adc_adc_slave_read;                        // mm_interconnect_0:adc_adc_slave_read -> adc:read
	wire         mm_interconnect_0_adc_adc_slave_write;                       // mm_interconnect_0:adc_adc_slave_write -> adc:write
	wire  [31:0] mm_interconnect_0_adc_adc_slave_writedata;                   // mm_interconnect_0:adc_adc_slave_writedata -> adc:writedata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_1_control_slave_readdata;       // sysid_qsys_1:readdata -> mm_interconnect_0:sysid_qsys_1_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_1_control_slave_address;        // mm_interconnect_0:sysid_qsys_1_control_slave_address -> sysid_qsys_1:address
	wire  [31:0] mm_interconnect_0_nios_1_debug_mem_slave_readdata;           // nios_1:debug_mem_slave_readdata -> mm_interconnect_0:nios_1_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_1_debug_mem_slave_waitrequest;        // nios_1:debug_mem_slave_waitrequest -> mm_interconnect_0:nios_1_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_1_debug_mem_slave_debugaccess;        // mm_interconnect_0:nios_1_debug_mem_slave_debugaccess -> nios_1:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_1_debug_mem_slave_address;            // mm_interconnect_0:nios_1_debug_mem_slave_address -> nios_1:debug_mem_slave_address
	wire         mm_interconnect_0_nios_1_debug_mem_slave_read;               // mm_interconnect_0:nios_1_debug_mem_slave_read -> nios_1:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_1_debug_mem_slave_byteenable;         // mm_interconnect_0:nios_1_debug_mem_slave_byteenable -> nios_1:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_1_debug_mem_slave_write;              // mm_interconnect_0:nios_1_debug_mem_slave_write -> nios_1:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_1_debug_mem_slave_writedata;          // mm_interconnect_0:nios_1_debug_mem_slave_writedata -> nios_1:debug_mem_slave_writedata
	wire         mm_interconnect_0_flash_epcs_control_port_chipselect;        // mm_interconnect_0:flash_epcs_control_port_chipselect -> flash:chipselect
	wire  [31:0] mm_interconnect_0_flash_epcs_control_port_readdata;          // flash:readdata -> mm_interconnect_0:flash_epcs_control_port_readdata
	wire   [8:0] mm_interconnect_0_flash_epcs_control_port_address;           // mm_interconnect_0:flash_epcs_control_port_address -> flash:address
	wire         mm_interconnect_0_flash_epcs_control_port_read;              // mm_interconnect_0:flash_epcs_control_port_read -> flash:read_n
	wire         mm_interconnect_0_flash_epcs_control_port_write;             // mm_interconnect_0:flash_epcs_control_port_write -> flash:write_n
	wire  [31:0] mm_interconnect_0_flash_epcs_control_port_writedata;         // mm_interconnect_0:flash_epcs_control_port_writedata -> flash:writedata
	wire  [31:0] mm_interconnect_0_altpll_pll_slave_readdata;                 // altpll:readdata -> mm_interconnect_0:altpll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_pll_slave_address;                  // mm_interconnect_0:altpll_pll_slave_address -> altpll:address
	wire         mm_interconnect_0_altpll_pll_slave_read;                     // mm_interconnect_0:altpll_pll_slave_read -> altpll:read
	wire         mm_interconnect_0_altpll_pll_slave_write;                    // mm_interconnect_0:altpll_pll_slave_write -> altpll:write
	wire  [31:0] mm_interconnect_0_altpll_pll_slave_writedata;                // mm_interconnect_0:altpll_pll_slave_writedata -> altpll:writedata
	wire         mm_interconnect_0_led_s1_chipselect;                         // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                           // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;                            // mm_interconnect_0:led_s1_address -> led:address
	wire         mm_interconnect_0_led_s1_write;                              // mm_interconnect_0:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                          // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                       // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                         // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                      // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                          // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                             // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                       // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                    // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                            // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                        // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_uart_s1_chipselect;                        // mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                          // uart:readdata -> mm_interconnect_0:uart_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                           // mm_interconnect_0:uart_s1_address -> uart:address
	wire         mm_interconnect_0_uart_s1_read;                              // mm_interconnect_0:uart_s1_read -> uart:read_n
	wire         mm_interconnect_0_uart_s1_begintransfer;                     // mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	wire         mm_interconnect_0_uart_s1_write;                             // mm_interconnect_0:uart_s1_write -> uart:write_n
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;                         // mm_interconnect_0:uart_s1_writedata -> uart:writedata
	wire         mm_interconnect_0_onchip_1_s1_chipselect;                    // mm_interconnect_0:onchip_1_s1_chipselect -> onchip_1:chipselect
	wire  [31:0] mm_interconnect_0_onchip_1_s1_readdata;                      // onchip_1:readdata -> mm_interconnect_0:onchip_1_s1_readdata
	wire  [11:0] mm_interconnect_0_onchip_1_s1_address;                       // mm_interconnect_0:onchip_1_s1_address -> onchip_1:address
	wire   [3:0] mm_interconnect_0_onchip_1_s1_byteenable;                    // mm_interconnect_0:onchip_1_s1_byteenable -> onchip_1:byteenable
	wire         mm_interconnect_0_onchip_1_s1_write;                         // mm_interconnect_0:onchip_1_s1_write -> onchip_1:write
	wire  [31:0] mm_interconnect_0_onchip_1_s1_writedata;                     // mm_interconnect_0:onchip_1_s1_writedata -> onchip_1:writedata
	wire         mm_interconnect_0_onchip_1_s1_clken;                         // mm_interconnect_0:onchip_1_s1_clken -> onchip_1:clken
	wire         mm_interconnect_0_spi_0_spi_control_port_chipselect;         // mm_interconnect_0:spi_0_spi_control_port_chipselect -> spi_0:spi_select
	wire  [31:0] mm_interconnect_0_spi_0_spi_control_port_readdata;           // spi_0:data_to_cpu -> mm_interconnect_0:spi_0_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_0_spi_control_port_address;            // mm_interconnect_0:spi_0_spi_control_port_address -> spi_0:mem_addr
	wire         mm_interconnect_0_spi_0_spi_control_port_read;               // mm_interconnect_0:spi_0_spi_control_port_read -> spi_0:read_n
	wire         mm_interconnect_0_spi_0_spi_control_port_write;              // mm_interconnect_0:spi_0_spi_control_port_write -> spi_0:write_n
	wire  [31:0] mm_interconnect_0_spi_0_spi_control_port_writedata;          // mm_interconnect_0:spi_0_spi_control_port_writedata -> spi_0:data_from_cpu
	wire  [31:0] mm_interconnect_0_nios_2_debug_mem_slave_readdata;           // nios_2:debug_mem_slave_readdata -> mm_interconnect_0:nios_2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_2_debug_mem_slave_waitrequest;        // nios_2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios_2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_2_debug_mem_slave_debugaccess;        // mm_interconnect_0:nios_2_debug_mem_slave_debugaccess -> nios_2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_2_debug_mem_slave_address;            // mm_interconnect_0:nios_2_debug_mem_slave_address -> nios_2:debug_mem_slave_address
	wire         mm_interconnect_0_nios_2_debug_mem_slave_read;               // mm_interconnect_0:nios_2_debug_mem_slave_read -> nios_2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_2_debug_mem_slave_byteenable;         // mm_interconnect_0:nios_2_debug_mem_slave_byteenable -> nios_2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_2_debug_mem_slave_write;              // mm_interconnect_0:nios_2_debug_mem_slave_write -> nios_2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_2_debug_mem_slave_writedata;          // mm_interconnect_0:nios_2_debug_mem_slave_writedata -> nios_2:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_2_s1_chipselect;                    // mm_interconnect_0:onchip_2_s1_chipselect -> onchip_2:chipselect
	wire  [31:0] mm_interconnect_0_onchip_2_s1_readdata;                      // onchip_2:readdata -> mm_interconnect_0:onchip_2_s1_readdata
	wire  [11:0] mm_interconnect_0_onchip_2_s1_address;                       // mm_interconnect_0:onchip_2_s1_address -> onchip_2:address
	wire   [3:0] mm_interconnect_0_onchip_2_s1_byteenable;                    // mm_interconnect_0:onchip_2_s1_byteenable -> onchip_2:byteenable
	wire         mm_interconnect_0_onchip_2_s1_write;                         // mm_interconnect_0:onchip_2_s1_write -> onchip_2:write
	wire  [31:0] mm_interconnect_0_onchip_2_s1_writedata;                     // mm_interconnect_0:onchip_2_s1_writedata -> onchip_2:writedata
	wire         mm_interconnect_0_onchip_2_s1_clken;                         // mm_interconnect_0:onchip_2_s1_clken -> onchip_2:clken
	wire         irq_mapper_receiver1_irq;                                    // uart:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios_1_irq_irq;                                              // irq_mapper:sender_irq -> nios_1:irq
	wire  [31:0] nios_2_irq_irq;                                              // irq_mapper_001:sender_irq -> nios_2:irq
	wire         irq_mapper_receiver2_irq;                                    // flash:irq -> [irq_mapper:receiver2_irq, irq_mapper_001:receiver1_irq]
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> [irq_mapper:receiver0_irq, irq_mapper_001:receiver0_irq]
	wire         irq_mapper_receiver3_irq;                                    // spi_0:irq -> [irq_mapper:receiver3_irq, irq_mapper_001:receiver2_irq]
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [adc:reset, flash:reset_n, jtag_uart_0:rst_n, mm_interconnect_0:adc_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sdram:reset_n, spi_0:reset_n, sysid_qsys_1:reset_n, uart:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [flash:reset_req, rst_translator:reset_req_in]
	wire         nios_1_debug_reset_request_reset;                            // nios_1:debug_reset_request -> [rst_controller:reset_in1, rst_controller_002:reset_in1]
	wire         nios_2_debug_reset_request_reset;                            // nios_2:debug_reset_request -> [rst_controller:reset_in2, rst_controller_003:reset_in1]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [altpll:reset, mm_interconnect_0:altpll_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;                          // rst_controller_002:reset_out -> [irq_mapper:reset, led:reset_n, mm_interconnect_0:nios_1_reset_reset_bridge_in_reset_reset, nios_1:reset_n, onchip_1:reset, rst_translator_001:in_reset]
	wire         rst_controller_002_reset_out_reset_req;                      // rst_controller_002:reset_req -> [nios_1:reset_req, onchip_1:reset_req, rst_translator_001:reset_req_in]
	wire         rst_controller_003_reset_out_reset;                          // rst_controller_003:reset_out -> [irq_mapper_001:reset, mm_interconnect_0:nios_2_reset_reset_bridge_in_reset_reset, nios_2:reset_n, onchip_2:reset]
	wire         rst_controller_003_reset_out_reset_req;                      // rst_controller_003:reset_req -> [nios_2:reset_req, onchip_2:reset_req, rst_translator_002:reset_req_in]

	helen_adc #(
		.board          ("DE0-Nano"),
		.board_rev      ("Autodetect"),
		.tsclk          (31),
		.numch          (8),
		.max10pllmultby (1),
		.max10plldivby  (1)
	) adc (
		.clock       (altpll_c0_clk),                               //                clk.clk
		.reset       (rst_controller_reset_out_reset),              //              reset.reset
		.write       (mm_interconnect_0_adc_adc_slave_write),       //          adc_slave.write
		.readdata    (mm_interconnect_0_adc_adc_slave_readdata),    //                   .readdata
		.writedata   (mm_interconnect_0_adc_adc_slave_writedata),   //                   .writedata
		.address     (mm_interconnect_0_adc_adc_slave_address),     //                   .address
		.waitrequest (mm_interconnect_0_adc_adc_slave_waitrequest), //                   .waitrequest
		.read        (mm_interconnect_0_adc_adc_slave_read),        //                   .read
		.adc_sclk    (adc_sclk),                                    // external_interface.export
		.adc_cs_n    (adc_cs_n),                                    //                   .export
		.adc_dout    (adc_dout),                                    //                   .export
		.adc_din     (adc_din)                                      //                   .export
	);

	helen_altpll altpll (
		.clk                (clk_clk),                                      //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),           // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_c0_clk),                                //                    c0.clk
		.c1                 (altpll_sdram_clk),                             //                    c1.clk
		.areset             (altpll_areset_conduit_export),                 //        areset_conduit.export
		.locked             (altpll_locked_conduit_export),                 //        locked_conduit.export
		.scandone           (),                                             //           (terminated)
		.scandataout        (),                                             //           (terminated)
		.phasedone          (),                                             //           (terminated)
		.phasecounterselect (4'b0000),                                      //           (terminated)
		.phaseupdown        (1'b0),                                         //           (terminated)
		.phasestep          (1'b0),                                         //           (terminated)
		.scanclk            (1'b0),                                         //           (terminated)
		.scanclkena         (1'b0),                                         //           (terminated)
		.scandata           (1'b0),                                         //           (terminated)
		.configupdate       (1'b0)                                          //           (terminated)
	);

	helen_flash flash (
		.clk        (altpll_c0_clk),                                        //               clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.reset_req  (rst_controller_reset_out_reset_req),                   //                  .reset_req
		.address    (mm_interconnect_0_flash_epcs_control_port_address),    // epcs_control_port.address
		.chipselect (mm_interconnect_0_flash_epcs_control_port_chipselect), //                  .chipselect
		.read_n     (~mm_interconnect_0_flash_epcs_control_port_read),      //                  .read_n
		.readdata   (mm_interconnect_0_flash_epcs_control_port_readdata),   //                  .readdata
		.write_n    (~mm_interconnect_0_flash_epcs_control_port_write),     //                  .write_n
		.writedata  (mm_interconnect_0_flash_epcs_control_port_writedata),  //                  .writedata
		.irq        (irq_mapper_receiver2_irq),                             //               irq.irq
		.dclk       (flash_dclk),                                           //          external.export
		.sce        (flash_sce),                                            //                  .export
		.sdo        (flash_sdo),                                            //                  .export
		.data0      (flash_data0)                                           //                  .export
	);

	helen_jtag_uart_0 jtag_uart_0 (
		.clk            (altpll_c0_clk),                                               //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	helen_led led (
		.clk        (altpll_c0_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (ledg_export)                          // external_connection.export
	);

	helen_nios_1 nios_1 (
		.clk                                 (altpll_c0_clk),                                        //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),                  //                     reset.reset_n
		.reset_req                           (rst_controller_002_reset_out_reset_req),               //                          .reset_req
		.d_address                           (nios_1_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_1_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_1_data_master_read),                              //                          .read
		.d_readdata                          (nios_1_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_1_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_1_data_master_write),                             //                          .write
		.d_writedata                         (nios_1_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios_1_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_1_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_1_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_1_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_1_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios_1_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios_1_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_1_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_1_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_1_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_1_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_1_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_1_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_1_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_1_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                      // custom_instruction_master.readra
	);

	helen_nios_2 nios_2 (
		.clk                                 (altpll_c0_clk),                                        //                       clk.clk
		.reset_n                             (~rst_controller_003_reset_out_reset),                  //                     reset.reset_n
		.reset_req                           (rst_controller_003_reset_out_reset_req),               //                          .reset_req
		.d_address                           (nios_2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_2_data_master_read),                              //                          .read
		.d_readdata                          (nios_2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_2_data_master_write),                             //                          .write
		.d_writedata                         (nios_2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios_2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_2_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios_2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios_2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                      // custom_instruction_master.readra
	);

	helen_onchip_1 onchip_1 (
		.clk        (altpll_c0_clk),                            //   clk1.clk
		.address    (mm_interconnect_0_onchip_1_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_1_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_1_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_1_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_1_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_1_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_1_s1_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),       // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req),   //       .reset_req
		.freeze     (1'b0)                                      // (terminated)
	);

	helen_onchip_2 onchip_2 (
		.clk        (altpll_c0_clk),                            //   clk1.clk
		.address    (mm_interconnect_0_onchip_2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_003_reset_out_reset),       // reset1.reset
		.reset_req  (rst_controller_003_reset_out_reset_req),   //       .reset_req
		.freeze     (1'b0)                                      // (terminated)
	);

	helen_sdram sdram (
		.clk            (altpll_c0_clk),                            //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	helen_spi_0 spi_0 (
		.clk           (altpll_c0_clk),                                       //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                     //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_0_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_0_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_0_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_0_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_0_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_0_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver3_irq),                            //              irq.irq
		.MISO          (spi_MISO),                                            //         external.export
		.MOSI          (spi_MOSI),                                            //                 .export
		.SCLK          (spi_SCLK),                                            //                 .export
		.SS_n          (spi_SS_n)                                             //                 .export
	);

	helen_sysid_qsys_1 sysid_qsys_1 (
		.clock    (altpll_c0_clk),                                         //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_1_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_1_control_slave_address)   //              .address
	);

	helen_uart uart (
		.clk           (altpll_c0_clk),                           //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.rxd           (uart_rxd),                                // external_connection.export
		.txd           (uart_txd),                                //                    .export
		.irq           (irq_mapper_receiver1_irq)                 //                 irq.irq
	);

	helen_mm_interconnect_0 mm_interconnect_0 (
		.altpll_c0_clk                                            (altpll_c0_clk),                                               //                                          altpll_c0.clk
		.clk_clk_clk                                              (clk_clk),                                                     //                                            clk_clk.clk
		.adc_reset_reset_bridge_in_reset_reset                    (rst_controller_reset_out_reset),                              //                    adc_reset_reset_bridge_in_reset.reset
		.altpll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // altpll_inclk_interface_reset_reset_bridge_in_reset.reset
		.nios_1_reset_reset_bridge_in_reset_reset                 (rst_controller_002_reset_out_reset),                          //                 nios_1_reset_reset_bridge_in_reset.reset
		.nios_2_reset_reset_bridge_in_reset_reset                 (rst_controller_003_reset_out_reset),                          //                 nios_2_reset_reset_bridge_in_reset.reset
		.nios_1_data_master_address                               (nios_1_data_master_address),                                  //                                 nios_1_data_master.address
		.nios_1_data_master_waitrequest                           (nios_1_data_master_waitrequest),                              //                                                   .waitrequest
		.nios_1_data_master_byteenable                            (nios_1_data_master_byteenable),                               //                                                   .byteenable
		.nios_1_data_master_read                                  (nios_1_data_master_read),                                     //                                                   .read
		.nios_1_data_master_readdata                              (nios_1_data_master_readdata),                                 //                                                   .readdata
		.nios_1_data_master_write                                 (nios_1_data_master_write),                                    //                                                   .write
		.nios_1_data_master_writedata                             (nios_1_data_master_writedata),                                //                                                   .writedata
		.nios_1_data_master_debugaccess                           (nios_1_data_master_debugaccess),                              //                                                   .debugaccess
		.nios_1_instruction_master_address                        (nios_1_instruction_master_address),                           //                          nios_1_instruction_master.address
		.nios_1_instruction_master_waitrequest                    (nios_1_instruction_master_waitrequest),                       //                                                   .waitrequest
		.nios_1_instruction_master_read                           (nios_1_instruction_master_read),                              //                                                   .read
		.nios_1_instruction_master_readdata                       (nios_1_instruction_master_readdata),                          //                                                   .readdata
		.nios_2_data_master_address                               (nios_2_data_master_address),                                  //                                 nios_2_data_master.address
		.nios_2_data_master_waitrequest                           (nios_2_data_master_waitrequest),                              //                                                   .waitrequest
		.nios_2_data_master_byteenable                            (nios_2_data_master_byteenable),                               //                                                   .byteenable
		.nios_2_data_master_read                                  (nios_2_data_master_read),                                     //                                                   .read
		.nios_2_data_master_readdata                              (nios_2_data_master_readdata),                                 //                                                   .readdata
		.nios_2_data_master_write                                 (nios_2_data_master_write),                                    //                                                   .write
		.nios_2_data_master_writedata                             (nios_2_data_master_writedata),                                //                                                   .writedata
		.nios_2_data_master_debugaccess                           (nios_2_data_master_debugaccess),                              //                                                   .debugaccess
		.nios_2_instruction_master_address                        (nios_2_instruction_master_address),                           //                          nios_2_instruction_master.address
		.nios_2_instruction_master_waitrequest                    (nios_2_instruction_master_waitrequest),                       //                                                   .waitrequest
		.nios_2_instruction_master_read                           (nios_2_instruction_master_read),                              //                                                   .read
		.nios_2_instruction_master_readdata                       (nios_2_instruction_master_readdata),                          //                                                   .readdata
		.adc_adc_slave_address                                    (mm_interconnect_0_adc_adc_slave_address),                     //                                      adc_adc_slave.address
		.adc_adc_slave_write                                      (mm_interconnect_0_adc_adc_slave_write),                       //                                                   .write
		.adc_adc_slave_read                                       (mm_interconnect_0_adc_adc_slave_read),                        //                                                   .read
		.adc_adc_slave_readdata                                   (mm_interconnect_0_adc_adc_slave_readdata),                    //                                                   .readdata
		.adc_adc_slave_writedata                                  (mm_interconnect_0_adc_adc_slave_writedata),                   //                                                   .writedata
		.adc_adc_slave_waitrequest                                (mm_interconnect_0_adc_adc_slave_waitrequest),                 //                                                   .waitrequest
		.altpll_pll_slave_address                                 (mm_interconnect_0_altpll_pll_slave_address),                  //                                   altpll_pll_slave.address
		.altpll_pll_slave_write                                   (mm_interconnect_0_altpll_pll_slave_write),                    //                                                   .write
		.altpll_pll_slave_read                                    (mm_interconnect_0_altpll_pll_slave_read),                     //                                                   .read
		.altpll_pll_slave_readdata                                (mm_interconnect_0_altpll_pll_slave_readdata),                 //                                                   .readdata
		.altpll_pll_slave_writedata                               (mm_interconnect_0_altpll_pll_slave_writedata),                //                                                   .writedata
		.flash_epcs_control_port_address                          (mm_interconnect_0_flash_epcs_control_port_address),           //                            flash_epcs_control_port.address
		.flash_epcs_control_port_write                            (mm_interconnect_0_flash_epcs_control_port_write),             //                                                   .write
		.flash_epcs_control_port_read                             (mm_interconnect_0_flash_epcs_control_port_read),              //                                                   .read
		.flash_epcs_control_port_readdata                         (mm_interconnect_0_flash_epcs_control_port_readdata),          //                                                   .readdata
		.flash_epcs_control_port_writedata                        (mm_interconnect_0_flash_epcs_control_port_writedata),         //                                                   .writedata
		.flash_epcs_control_port_chipselect                       (mm_interconnect_0_flash_epcs_control_port_chipselect),        //                                                   .chipselect
		.jtag_uart_0_avalon_jtag_slave_address                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                      jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                                   .write
		.jtag_uart_0_avalon_jtag_slave_read                       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                                   .read
		.jtag_uart_0_avalon_jtag_slave_readdata                   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                                   .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                                   .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                                   .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                 (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                                   .chipselect
		.led_s1_address                                           (mm_interconnect_0_led_s1_address),                            //                                             led_s1.address
		.led_s1_write                                             (mm_interconnect_0_led_s1_write),                              //                                                   .write
		.led_s1_readdata                                          (mm_interconnect_0_led_s1_readdata),                           //                                                   .readdata
		.led_s1_writedata                                         (mm_interconnect_0_led_s1_writedata),                          //                                                   .writedata
		.led_s1_chipselect                                        (mm_interconnect_0_led_s1_chipselect),                         //                                                   .chipselect
		.nios_1_debug_mem_slave_address                           (mm_interconnect_0_nios_1_debug_mem_slave_address),            //                             nios_1_debug_mem_slave.address
		.nios_1_debug_mem_slave_write                             (mm_interconnect_0_nios_1_debug_mem_slave_write),              //                                                   .write
		.nios_1_debug_mem_slave_read                              (mm_interconnect_0_nios_1_debug_mem_slave_read),               //                                                   .read
		.nios_1_debug_mem_slave_readdata                          (mm_interconnect_0_nios_1_debug_mem_slave_readdata),           //                                                   .readdata
		.nios_1_debug_mem_slave_writedata                         (mm_interconnect_0_nios_1_debug_mem_slave_writedata),          //                                                   .writedata
		.nios_1_debug_mem_slave_byteenable                        (mm_interconnect_0_nios_1_debug_mem_slave_byteenable),         //                                                   .byteenable
		.nios_1_debug_mem_slave_waitrequest                       (mm_interconnect_0_nios_1_debug_mem_slave_waitrequest),        //                                                   .waitrequest
		.nios_1_debug_mem_slave_debugaccess                       (mm_interconnect_0_nios_1_debug_mem_slave_debugaccess),        //                                                   .debugaccess
		.nios_2_debug_mem_slave_address                           (mm_interconnect_0_nios_2_debug_mem_slave_address),            //                             nios_2_debug_mem_slave.address
		.nios_2_debug_mem_slave_write                             (mm_interconnect_0_nios_2_debug_mem_slave_write),              //                                                   .write
		.nios_2_debug_mem_slave_read                              (mm_interconnect_0_nios_2_debug_mem_slave_read),               //                                                   .read
		.nios_2_debug_mem_slave_readdata                          (mm_interconnect_0_nios_2_debug_mem_slave_readdata),           //                                                   .readdata
		.nios_2_debug_mem_slave_writedata                         (mm_interconnect_0_nios_2_debug_mem_slave_writedata),          //                                                   .writedata
		.nios_2_debug_mem_slave_byteenable                        (mm_interconnect_0_nios_2_debug_mem_slave_byteenable),         //                                                   .byteenable
		.nios_2_debug_mem_slave_waitrequest                       (mm_interconnect_0_nios_2_debug_mem_slave_waitrequest),        //                                                   .waitrequest
		.nios_2_debug_mem_slave_debugaccess                       (mm_interconnect_0_nios_2_debug_mem_slave_debugaccess),        //                                                   .debugaccess
		.onchip_1_s1_address                                      (mm_interconnect_0_onchip_1_s1_address),                       //                                        onchip_1_s1.address
		.onchip_1_s1_write                                        (mm_interconnect_0_onchip_1_s1_write),                         //                                                   .write
		.onchip_1_s1_readdata                                     (mm_interconnect_0_onchip_1_s1_readdata),                      //                                                   .readdata
		.onchip_1_s1_writedata                                    (mm_interconnect_0_onchip_1_s1_writedata),                     //                                                   .writedata
		.onchip_1_s1_byteenable                                   (mm_interconnect_0_onchip_1_s1_byteenable),                    //                                                   .byteenable
		.onchip_1_s1_chipselect                                   (mm_interconnect_0_onchip_1_s1_chipselect),                    //                                                   .chipselect
		.onchip_1_s1_clken                                        (mm_interconnect_0_onchip_1_s1_clken),                         //                                                   .clken
		.onchip_2_s1_address                                      (mm_interconnect_0_onchip_2_s1_address),                       //                                        onchip_2_s1.address
		.onchip_2_s1_write                                        (mm_interconnect_0_onchip_2_s1_write),                         //                                                   .write
		.onchip_2_s1_readdata                                     (mm_interconnect_0_onchip_2_s1_readdata),                      //                                                   .readdata
		.onchip_2_s1_writedata                                    (mm_interconnect_0_onchip_2_s1_writedata),                     //                                                   .writedata
		.onchip_2_s1_byteenable                                   (mm_interconnect_0_onchip_2_s1_byteenable),                    //                                                   .byteenable
		.onchip_2_s1_chipselect                                   (mm_interconnect_0_onchip_2_s1_chipselect),                    //                                                   .chipselect
		.onchip_2_s1_clken                                        (mm_interconnect_0_onchip_2_s1_clken),                         //                                                   .clken
		.sdram_s1_address                                         (mm_interconnect_0_sdram_s1_address),                          //                                           sdram_s1.address
		.sdram_s1_write                                           (mm_interconnect_0_sdram_s1_write),                            //                                                   .write
		.sdram_s1_read                                            (mm_interconnect_0_sdram_s1_read),                             //                                                   .read
		.sdram_s1_readdata                                        (mm_interconnect_0_sdram_s1_readdata),                         //                                                   .readdata
		.sdram_s1_writedata                                       (mm_interconnect_0_sdram_s1_writedata),                        //                                                   .writedata
		.sdram_s1_byteenable                                      (mm_interconnect_0_sdram_s1_byteenable),                       //                                                   .byteenable
		.sdram_s1_readdatavalid                                   (mm_interconnect_0_sdram_s1_readdatavalid),                    //                                                   .readdatavalid
		.sdram_s1_waitrequest                                     (mm_interconnect_0_sdram_s1_waitrequest),                      //                                                   .waitrequest
		.sdram_s1_chipselect                                      (mm_interconnect_0_sdram_s1_chipselect),                       //                                                   .chipselect
		.spi_0_spi_control_port_address                           (mm_interconnect_0_spi_0_spi_control_port_address),            //                             spi_0_spi_control_port.address
		.spi_0_spi_control_port_write                             (mm_interconnect_0_spi_0_spi_control_port_write),              //                                                   .write
		.spi_0_spi_control_port_read                              (mm_interconnect_0_spi_0_spi_control_port_read),               //                                                   .read
		.spi_0_spi_control_port_readdata                          (mm_interconnect_0_spi_0_spi_control_port_readdata),           //                                                   .readdata
		.spi_0_spi_control_port_writedata                         (mm_interconnect_0_spi_0_spi_control_port_writedata),          //                                                   .writedata
		.spi_0_spi_control_port_chipselect                        (mm_interconnect_0_spi_0_spi_control_port_chipselect),         //                                                   .chipselect
		.sysid_qsys_1_control_slave_address                       (mm_interconnect_0_sysid_qsys_1_control_slave_address),        //                         sysid_qsys_1_control_slave.address
		.sysid_qsys_1_control_slave_readdata                      (mm_interconnect_0_sysid_qsys_1_control_slave_readdata),       //                                                   .readdata
		.uart_s1_address                                          (mm_interconnect_0_uart_s1_address),                           //                                            uart_s1.address
		.uart_s1_write                                            (mm_interconnect_0_uart_s1_write),                             //                                                   .write
		.uart_s1_read                                             (mm_interconnect_0_uart_s1_read),                              //                                                   .read
		.uart_s1_readdata                                         (mm_interconnect_0_uart_s1_readdata),                          //                                                   .readdata
		.uart_s1_writedata                                        (mm_interconnect_0_uart_s1_writedata),                         //                                                   .writedata
		.uart_s1_begintransfer                                    (mm_interconnect_0_uart_s1_begintransfer),                     //                                                   .begintransfer
		.uart_s1_chipselect                                       (mm_interconnect_0_uart_s1_chipselect)                         //                                                   .chipselect
	);

	helen_irq_mapper irq_mapper (
		.clk           (altpll_c0_clk),                      //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (nios_1_irq_irq)                      //    sender.irq
	);

	helen_irq_mapper_001 irq_mapper_001 (
		.clk           (altpll_c0_clk),                      //       clk.clk
		.reset         (rst_controller_003_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver2_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver3_irq),           // receiver2.irq
		.sender_irq    (nios_2_irq_irq)                      //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios_1_debug_reset_request_reset),   // reset_in1.reset
		.reset_in2      (nios_2_debug_reset_request_reset),   // reset_in2.reset
		.clk            (altpll_c0_clk),                      //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios_1_debug_reset_request_reset),       // reset_in1.reset
		.clk            (altpll_c0_clk),                          //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios_2_debug_reset_request_reset),       // reset_in1.reset
		.clk            (altpll_c0_clk),                          //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_003_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
