module led(
	LEDG
);

output [7:0] LEDG;

assign LEDG[1] = 1'b1;
endmodule